`ifndef LIB_TESTBENCH_SVH
`define LIB_TESTBENCH_SVH

`timescale 1ns/100ps

`define TIMESPEC      1e9
`define PERIOD_CALC(x) (`TIMESPEC/x)

`define LIB_CLK_GEN(name, period) logic name = 1'b0; always#(`PERIOD_CALC(period)/2.0) name++;
`define LIB_RST_GEN(rst_name, clk, delay_cycles) logic rst_name; initial begin rst_name = 1'b0; repeat(delay_cycles) @(posedge clk); rst_name = 1'b1; end
`define LIB_DUT_DRIVE_AXI4_STREAM_REAL(valid_name, last_name, data_name, data_width, clk, rst_n, data_queue) logic valid_name; logic last_name; logic signed [data_width-1:0] data_name; initial begin valid_name = 1'b0; last_name = 1'b0; data_name = '0; wait (rst_n === 1'b1); if (data_queue.size() > 0) begin for (int i = 0; i < data_queue.size(); i++) begin @(posedge clk); valid_name <= 1'b1; data_name  <= data_queue[i]; if (i == data_queue.size() - 1) begin last_name <= 1'b1; end end @(posedge clk); valid_name <= 1'b0; last_name  <= 1'b0; data_name  <= '0; end end
`define LIB_DUT_DRIVE_AXI4_STREAM_REAL_VERIFY(valid_name, last_name, data_name, data_width, clk, rst_n, data_queue) logic valid_name; logic last_name; logic signed [data_width-1:0] data_name; initial begin valid_name = 1'b0; last_name = 1'b0; data_name = '0; wait (rst_n === 1'b1); if (data_queue.size() > 0) begin int data_idx = 0; while (data_idx < data_queue.size()) begin @(posedge clk); if ($urandom_range(1, 10) > 5) begin valid_name <= 1'b1; data_name  <= data_queue[data_idx]; if (data_idx == data_queue.size() - 1) begin last_name <= 1'b1; end data_idx++; end else begin valid_name <= 1'b0; last_name  <= 1'b0; data_name  <= '0; end end @(posedge clk); valid_name <= 1'b0; last_name  <= 1'b0; data_name  <= '0; end end
`define LIB_DUT_DRIVE_AXI4_STREAM_COMPLEX(valid_name, last_name, data_name_real, data_name_imag, data_width, clk, rst_n, data_queue_real, data_queue_imag) logic valid_name; logic last_name; logic signed [data_width-1:0] data_name_real; logic signed [data_width-1:0] data_name_imag; initial begin valid_name = 1'b0; last_name = 1'b0; data_name_real = '0; data_name_imag = '0; wait (rst_n === 1'b1); assert (data_queue_real.size() == data_queue_imag.size()) else $fatal(1, "Complex AXI Stream queues must have the same size."); if (data_queue_real.size() > 0) begin for (int i = 0; i < data_queue_real.size(); i++) begin @(posedge clk); valid_name <= 1'b1; data_name_real <= data_queue_real[i]; data_name_imag <= data_queue_imag[i]; if (i == data_queue_real.size() - 1) begin last_name <= 1'b1; end end @(posedge clk); valid_name <= 1'b0; last_name  <= 1'b0; data_name_real <= '0; data_name_imag <= '0; end end
`define LIB_DUT_DRIVE_AXI4_STREAM_COMPLEX_VERIFY(valid_name, last_name, data_name_real, data_name_imag, data_width, clk, rst_n, data_queue_real, data_queue_imag) logic valid_name; logic last_name; logic signed [data_width-1:0] data_name_real; logic signed [data_width-1:0] data_name_imag; initial begin valid_name = 1'b0; last_name = 1'b0; data_name_real = '0; data_name_imag = '0; wait (rst_n === 1'b1); assert (data_queue_real.size() == data_queue_imag.size()) else $fatal(1, "Complex AXI Stream queues must have the same size."); if (data_queue_real.size() > 0) begin int data_idx = 0; while (data_idx < data_queue_real.size()) begin @(posedge clk); if ($urandom_range(1, 10) > 5) begin valid_name <= 1'b1; data_name_real <= data_queue_real[data_idx]; data_name_imag <= data_queue_imag[data_idx]; if (data_idx == data_queue_real.size() - 1) begin last_name <= 1'b1; end data_idx++; end else begin valid_name <= 1'b0; last_name  <= 1'b0; data_name_real <= '0; data_name_imag <= '0; end end @(posedge clk); valid_name <= 1'b0; last_name  <= 1'b0; data_name_real <= '0; data_name_imag <= '0; end end
`define LIB_DUT_TEST_VECTOR_FILE_READ(file_path, queue_mem) int queue_mem[$] = {}; initial begin int fd; int temp_val; int ret; fd = $fopen(file_path, "r"); if (fd == 0) begin $display("ERROR: File could not be opened: %s", file_path); $finish; end forever begin ret = $fscanf(fd, "%d\n", temp_val); if (ret != 1) break; queue_mem.push_back(temp_val); end $fclose(fd); end
`define LIB_DUT_OUTPUT_TO_FILE(clk, rst_n, valid_signal, data_signal, last_signal, filepath) initial begin integer output_file; wait (rst_n === 1'b1); output_file = $fopen(filepath, "w"); if (output_file == 0) begin $display("ERROR: %s 파일을 열 수 없습니다.", filepath); $finish; end fork forever @(posedge clk) begin if (rst_n && valid_signal) begin $fdisplay(output_file, "%d", data_signal); end end begin wait (last_signal === 1'b1); repeat(200) @(posedge clk); $fclose(output_file); $display("시뮬레이션 결과 저장이 완료되었습니다. -> %s", filepath); end join end
`define LIB_COMPARE_WITH_GOLDEN_REAL(clk, rst_n, valid_signal, data_signal, last_signal, golden_filepath) initial begin int golden_queue[$] = {}; int dut_output_queue[$] = {}; integer golden_file; integer temp_val; integer ret; integer mismatches = 0; int compare_size; golden_file = $fopen(golden_filepath, "r"); if (golden_file == 0) begin $display("ERROR: Golden Reference 파일을 열 수 없습니다: %s", golden_filepath); $finish; end while ($fscanf(golden_file, "%d\n", temp_val) == 1) begin golden_queue.push_back(temp_val); end $fclose(golden_file); wait (rst_n === 1'b1); forever @(posedge clk) begin if (rst_n && valid_signal) begin dut_output_queue.push_back(data_signal); if (last_signal) begin break; end end end repeat(10) @(posedge clk); $display("--- Golden Reference 비교 시작 ---"); if (golden_queue.size() != dut_output_queue.size()) begin $display("ERROR: 출력 데이터 개수가 다릅니다. Golden: %0d, DUT: %0d", golden_queue.size(), dut_output_queue.size()); mismatches++; end compare_size = (golden_queue.size() < dut_output_queue.size()) ? golden_queue.size() : dut_output_queue.size(); for (int i = 0; i < compare_size; i++) begin if (golden_queue[i] != dut_output_queue[i]) begin $display("ERROR: 데이터 불일치 (인덱스 %0d). Golden: %d, DUT: %d", i, golden_queue[i], dut_output_queue[i]); mismatches++; end end if (mismatches == 0) begin $display("SUCCESS: 결과가 일치합니다! (총 %0d개 데이터)", dut_output_queue.size()); end else begin $display("FAILURE: 총 %0d개의 불일치가 발견되었습니다.", mismatches); end $display("------------------------------------"); $finish; end
`define LIB_COMPARE_WITH_GOLDEN_COMPLEX(clk, rst_n, valid_signal, data_signal_real, data_signal_imag, last_signal, golden_filepath_real, golden_filepath_imag) initial begin int golden_queue_real[$] = {}; int golden_queue_imag[$] = {}; int dut_output_queue_real[$] = {}; int dut_output_queue_imag[$] = {}; integer golden_file; integer temp_val; integer mismatches = 0; int compare_size; golden_file = $fopen(golden_filepath_real, "r"); if (golden_file == 0) begin $display("ERROR: Golden Real 파일을 열 수 없습니다: %s", golden_filepath_real); $finish; end while ($fscanf(golden_file, "%d\n", temp_val) == 1) begin golden_queue_real.push_back(temp_val); end $fclose(golden_file); golden_file = $fopen(golden_filepath_imag, "r"); if (golden_file == 0) begin $display("ERROR: Golden Imaginary 파일을 열 수 없습니다: %s", golden_filepath_imag); $finish; end while ($fscanf(golden_file, "%d\n", temp_val) == 1) begin golden_queue_imag.push_back(temp_val); end $fclose(golden_file); assert (golden_queue_real.size() == golden_queue_imag.size()) else $fatal(1, "실수부와 허수부 골든 파일의 데이터 개수가 다릅니다."); wait (rst_n === 1'b1); forever @(posedge clk) begin if (rst_n && valid_signal) begin dut_output_queue_real.push_back(data_signal_real); dut_output_queue_imag.push_back(data_signal_imag); if (last_signal) begin break; end end end repeat(10) @(posedge clk); $display("--- Golden Reference 비교 시작 (복소수) ---"); if (golden_queue_real.size() != dut_output_queue_real.size()) begin $display("ERROR: 출력 데이터 개수가 다릅니다. Golden: %0d, DUT: %0d", golden_queue_real.size(), dut_output_queue_real.size()); mismatches++; end compare_size = (golden_queue_real.size() < dut_output_queue_real.size()) ? golden_queue_real.size() : dut_output_queue_real.size(); for (int i = 0; i < compare_size; i++) begin if (golden_queue_real[i] != dut_output_queue_real[i]) begin $display("ERROR: [실수부] 데이터 불일치 (인덱스 %0d). Golden: %d, DUT: %d", i, golden_queue_real[i], dut_output_queue_real[i]); mismatches++; end if (golden_queue_imag[i] != dut_output_queue_imag[i]) begin $display("ERROR: [허수부] 데이터 불일치 (인덱스 %0d). Golden: %d, DUT: %d", i, golden_queue_imag[i], dut_output_queue_imag[i]); mismatches++; end end if (mismatches == 0) begin $display("SUCCESS: 결과가 일치합니다! (총 %0d개 복소수 데이터)", dut_output_queue_real.size()); end else begin $display("FAILURE: 총 %0d개의 불일치가 발견되었습니다.", mismatches); end $display("-------------------------------------------"); $finish; end

`endif // LIB_TESTBENCH_SVH
